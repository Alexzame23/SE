library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity image is
    port(
        clk_108mhz          : in  std_logic;
        reset_n             : in  std_logic;
        row, col            : in  std_logic_vector(15 downto 0);
        rout, gout, bout    : out std_logic_vector(3 downto 0);
         row_new_pixel: in  std_logic_vector(3 downto 0);
          col_new_pixel: in  std_logic_vector(3 downto 0);
              load_new_pixel      : in  std_logic;
            color_new_pixel     : in  std_logic_vector(11 downto 0));
end entity;

architecture arch of image is
--    type ram_type is array (0 to 65536-1) of std_logic_vector(11 downto 0);
      type ram_type is array (0 to 256-1) of std_logic_vector(11 downto 0);
    signal RAM : ram_type :=
    (
    "111100000000", "000000001111", "111100000000", "000000001111", "111100000000", "000000001111","111100000000","000000001111",
    "111100000000", "000000001111", "111100000000", "000000001111", "111100000000","000000001111","111100000000", "000000001111", 
    "000000001111", "111100000000", "000000001111", "111100000000", "000000001111","111100000000", "000000001111", "111100000000", 
    "000000001111", "111100000000", "000000001111", "111100000000","000000001111", "111100000000", "000000001111","111100000000",
    "111100000000", "000000001111","111100000000", "000000001111", "111100000000", "000000001111", "111100000000", "000000001111", 
    "111100000000","000000001111", "111100000000", "000000001111", "111100000000", "000000001111", "111100000000", "000000001111",
    "000000001111", "111100000000", "000000001111", "111100000000", "000000001111", "111100000000","000000001111","111100000000", 
    "000000001111", "111100000000", "000000001111", "111100000000", "000000001111","111100000000", "000000001111", "111100000000", 
    "111100000000", "000000001111", "111100000000","000000001111", "111100000000", "000000001111", "111100000000", "000000001111", 
    "111100000000", "000000001111","111100000000","000000001111", "111100000000", "000000001111", "111100000000", "000000001111", 
    "000000001111", "111100000000", "000000001111", "111100000000", "000000001111", "111100000000", "000000001111","111100000000",
    "000000001111", "111100000000", "000000001111", "111100000000", "000000001111", "111100000000","000000001111","111100000000", 
    "111100000000", "000000001111", "111100000000", "000000001111","111100000000", "000000001111", "111100000000", "000000001111",
    "111100000000", "000000001111", "111100000000","000000001111","111100000000", "000000001111", "111100000000", "000000001111", 
    "000000001111","111100000000", "000000001111", "111100000000", "000000001111", "111100000000", "000000001111", "111100000000",
    "000000001111","111100000000", "000000001111", "111100000000", "000000001111", "111100000000", "000000001111", "111100000000",
      "111100000000", "000000001111", "111100000000", "000000001111", "111100000000", "000000001111","111100000000","000000001111",
    "111100000000", "000000001111", "111100000000", "000000001111", "111100000000","000000001111","111100000000", "000000001111", 
    "000000001111", "111100000000", "000000001111", "111100000000", "000000001111","111100000000", "000000001111", "111100000000", 
    "000000001111", "111100000000", "000000001111", "111100000000","000000001111", "111100000000", "000000001111","111100000000",
    "111100000000", "000000001111","111100000000", "000000001111", "111100000000", "000000001111", "111100000000", "000000001111", 
    "111100000000","000000001111", "111100000000", "000000001111", "111100000000", "000000001111", "111100000000", "000000001111",
    "000000001111", "111100000000", "000000001111", "111100000000", "000000001111", "111100000000","000000001111","111100000000", 
    "000000001111", "111100000000", "000000001111", "111100000000", "000000001111","111100000000", "000000001111", "111100000000", 
    "111100000000", "000000001111", "111100000000","000000001111", "111100000000", "000000001111", "111100000000", "000000001111", 
    "111100000000", "000000001111","111100000000","000000001111", "111100000000", "000000001111", "111100000000", "000000001111", 
    "000000001111", "111100000000", "000000001111", "111100000000", "000000001111", "111100000000", "000000001111","111100000000",
    "000000001111", "111100000000", "000000001111", "111100000000", "000000001111", "111100000000","000000001111","111100000000", 
    "111100000000", "000000001111", "111100000000", "000000001111","111100000000", "000000001111", "111100000000", "000000001111",
    "111100000000", "000000001111", "111100000000","000000001111","111100000000", "000000001111", "111100000000", "000000001111", 
    "000000001111","111100000000", "000000001111", "111100000000", "000000001111", "111100000000", "000000001111", "111100000000",
    "000000001111","111100000000", "000000001111", "111100000000", "000000001111", "111100000000", "000000001111", "111100000000"
    
    );
    
--    signal row_and_col : std_logic_vector(15 downto 0);
        signal row_and_col, row_and_col_new_pixel : std_logic_vector(7 downto 0);
    
               
    
begin

 --   row_and_col <= row(7 downto 0) & col(7 downto 0);
    row_and_col <= row(7 downto 4) & col(7 downto 4);
       row_and_col_new_pixel <= row_new_pixel& col_new_pixel;
  
               process(clk_108mhz)
    begin
        if rising_edge(clk_108mhz) then
        if (load_new_pixel = '1' ) then 
            RAM(to_integer(unsigned(row_and_col_new_pixel)))(11 downto 8)<= color_new_pixel(11 downto 8);
             RAM(to_integer(unsigned(row_and_col_new_pixel)))( 7 downto 4)<= color_new_pixel(7 downto 4);
           RAM(to_integer(unsigned(row_and_col_new_pixel)))( 3 downto 0)<= color_new_pixel(3 downto 0);
           end if;
       end if;    
      end process;
    
   
    process(clk_108mhz)
    begin
        if rising_edge(clk_108mhz) then

 		if ( to_integer(unsigned(row(15 downto 8))) =0 and to_integer(unsigned(col(15 downto 8))) =0 ) then

                rout <= RAM(to_integer(unsigned(row_and_col)))(11 downto 8);
                gout <= RAM(to_integer(unsigned(row_and_col)))( 7 downto 4);
                bout <= RAM(to_integer(unsigned(row_and_col)))( 3 downto 0);
            else
                rout <= "0000";
                gout <= "0000";
                bout <= "0000";
            end if;
        end if;
    end process;
end arch;